`ifndef header_h
`define header_h

`define REG_S 32
`define REG_ADD_W 5
`define REG_DAT_W 32

// mem
`define MEM_ADD_W 32
`define MEM_DAT_W 8

`define INS_DAT_W 32

`endif

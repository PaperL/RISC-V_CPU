`ifndef header_h
`define header_h

// Memory
`define MEM_ADD_W 32
`define MEM_DAT_W 8

// Register
`define REG_S 32
`define REG_ADD_W 5
`define REG_DAT_W 32

// Instruction
`define INS_DAT_W 32
`define INS_OP_W 5

// Reordered Buffer
`define ROB_S 32
`define ROB_ADD_W 5

// Reservation Station
`define RS_S 32
`define RS_ADD_W 5

`endif

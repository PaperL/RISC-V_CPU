`include "header.vh" 
// ReOrdered Buffer Module
module rob (
           input wire clk,
           input wire rst,
           input wire en
       );

always @(posedge clk) begin
    if (rst) begin
        // todo
    end
    else if (en) begin
        // todo
    end
end

endmodule
